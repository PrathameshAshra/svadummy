<svg xmlns="http://www.w3.org/2000/svg" width="23.514" height="20" viewBox="0 0 23.514 20">
  <g id="Home_Icon" data-name="Home Icon" transform="translate(-5 -5.3)" style="isolation: isolate">
    <path id="Path_1" data-name="Path 1" d="M8.514,25.3V15.894H5.006c0-.006,0-.013-.006-.016Q10.872,10.588,16.751,5.3q5.877,5.291,11.764,10.588H24.987V25.3H19.105V18.249H14.4V25.3C12.436,25.3,10.478,25.3,8.514,25.3Z" fill="#fe7c7b"/>
  </g>
</svg>
